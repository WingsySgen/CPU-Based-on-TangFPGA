`define LEN 8
`define RSTEDGE negedge
`define _RSTEDGE posedge
