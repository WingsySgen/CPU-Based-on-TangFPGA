`define module_name SPI_MASTER_Top
