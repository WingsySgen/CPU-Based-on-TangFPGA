`define module_name UART_MASTER_Top
